module top;
  initial begin
    $display( "Yes I modified it! Hello World!" );
  end
endmodule
